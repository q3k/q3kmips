module qm_fetch(
    /// datapath
    // output instruction register
    output wire [31:0] do_IR,
    // output next pc
    output wire [31:0] do_NextPC
);

endmodule
